* nfet_vgid.spice — Vg–Id sweep for sky130_fd_pr__nfet_01v8 (WSL/Linux/Windows ngspice 35+)
* Requires environment variables:
*   export PDK_ROOT=/mnt/c/openlane/pdks
*   export PDK=sky130A
.lib "$::env(PDK_ROOT)/$::env(PDK)/libs.tech/ngspice/sky130.lib.spice" tt

.options TEMP=25
.options METHOD=trap

.param W=1u
.param L=0.15u
.param VDS_BIAS=0.8

* Node order: D G S B
Vd  D  0  {VDS_BIAS}
Vg  G  0  0
Vs  S  0  0
Vb  B  0  0

M1  D  G  S  B  sky130_fd_pr__nfet_01v8  w={W}  l={L}

* Sweep gate from 0 → 1.8 V (typical 01v8 device)
.dc Vg 0 1.8 0.01

.control
  set wr_singlescale
  set wr_vecnames
  run
  * Drain current flowing D→S (positive): minus branch of Vd source
  let Id = -i(Vd)
  wrdata nfet_vgid.csv v(g) Id
  quit
.endc

.end
