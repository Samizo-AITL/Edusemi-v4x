* FinFET 15nm model (BSIM-CMG level=54)
.model nfinfet nmos level=54
+ version = 4.8
+ nch = 1.5e-7
+ tox = 1.2e-9
+ finwidth = 8e-9
+ finheight = 35e-9
+ nfin = 3
+ vth0 = 0.42
+ u0 = 300
+ rdsw = 500
+ cgso = 1e-10
+ cgdo = 1e-10
+ cgbo = 5e-11
+ cf = 2e-15
+ rs = 200
+ rd = 200
+ vsat = 1.2e7
+ pdiblc1 = 1.5e-2
+ pdiblc2 = 1e-3
+ eta0 = 0.1
+ dvt0 = 0.15
+ dvt1 = 0.4
+ dvt2 = 0.05
+ delt = 0.01
+ lint = 1.5e-9
