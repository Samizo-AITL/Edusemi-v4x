* GAA 5nm model (BSIM-CMG level=54)
.model ngaa nmos level=54
+ version = 4.8
+ nch = 8e-8
+ tox = 0.8e-9
+ finwidth = 5e-9
+ finheight = 45e-9
+ nsheet = 3
+ sheets_sep = 5e-9
+ vth0 = 0.38
+ u0 = 250
+ rdsw = 600
+ cgso = 1e-10
+ cgdo = 1e-10
+ cgbo = 5e-11
+ cf = 2e-15
+ rs = 250
+ rd = 250
+ vsat = 1.5e7
+ pdiblc1 = 1.2e-2
+ pdiblc2 = 8e-4
+ eta0 = 0.08
+ dvt0 = 0.12
+ dvt1 = 0.35
+ dvt2 = 0.04
+ delt = 0.01
+ lint = 1.0e-9
