* CMOS Inverter using CFET Stack Model
.include cfet_stack_model.spice

Vdd vdd 0 DC 0.8
Vin in 0 DC 0.0

* Stacked PMOS (Top)
M1 out in vdd vdd pcfet L=10n W=120n

* Stacked NMOS (Bottom)
M2 out in 0 0 ncfet L=10n W=120n

.dc Vin 0 0.8 0.01
.print dc V(in) V(out)
.end
