* pfet_vgid.spice — Vg–Id sweep for sky130_fd_pr__pfet_01v8
* Requires environment variables:
*   export PDK_ROOT=/mnt/c/openlane/pdks
*   export PDK=sky130A
.lib "$::env(PDK_ROOT)/$::env(PDK)/libs.tech/ngspice/sky130.lib.spice" tt

.options TEMP=25
.options METHOD=trap

.param W=1u
.param L=0.15u
.param VDD=0.9

* Node order: D G S B
* PFET in p-well: Source/Bulk at VDD, Drain at 0
Vd  D  0   0
Vg  G  0   0
Vs  S  0   {VDD}
Vb  B  0   {VDD}

M1  D  G  S  B  sky130_fd_pr__pfet_01v8  w={W}  l={L}

* Sweep gate from 1.8 → 0 V (more conductive as gate lowers)
.dc Vg 1.8 0 -0.01

.control
  set wr_singlescale
  set wr_vecnames
  run
  * Use magnitude so output is positive
  let Id = abs(i(Vd))
  wrdata pfet_vgid.csv v(g) Id
  quit
.endc

.end
